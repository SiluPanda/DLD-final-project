--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:45:06 04/17/2018
-- Design Name:   
-- Module Name:   /home/encryptor/test_clock.vhd
-- Project Name:  encryptor
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: clockconverter
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY test_clock IS
END test_clock;
 
ARCHITECTURE behavior OF test_clock IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT clockconverter
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         n : IN  std_logic_vector(5 downto 0);
         b_c_out : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal n : std_logic_vector(5 downto 0) := (others => '0');

 	--Outputs
   signal b_c_out : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: clockconverter PORT MAP (
          clk => clk,
          reset => reset,
          n => n,
          b_c_out => b_c_out
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		reset <= '1';
      wait for 100 ns;
		reset <= '0';
		n <= "001000";

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
